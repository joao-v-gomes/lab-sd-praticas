library verilog;
use verilog.vl_types.all;
entity identificaIndvA_vlg_check_tst is
    port(
        A               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end identificaIndvA_vlg_check_tst;
