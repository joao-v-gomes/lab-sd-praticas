library verilog;
use verilog.vl_types.all;
entity identificaIndvA_vlg_vec_tst is
end identificaIndvA_vlg_vec_tst;
