library verilog;
use verilog.vl_types.all;
entity Cofre_vhdl_vlg_vec_tst is
end Cofre_vhdl_vlg_vec_tst;
