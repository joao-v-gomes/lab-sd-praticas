library verilog;
use verilog.vl_types.all;
entity identificaIndvA is
    port(
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        D4              : in     vl_logic;
        D5              : in     vl_logic;
        L1              : in     vl_logic;
        L2              : in     vl_logic;
        L3              : in     vl_logic;
        L4              : in     vl_logic;
        L5              : in     vl_logic;
        A               : out    vl_logic
    );
end identificaIndvA;
