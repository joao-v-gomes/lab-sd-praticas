library verilog;
use verilog.vl_types.all;
entity andGate_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end andGate_vlg_check_tst;
